LCD.v